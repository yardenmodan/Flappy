module Buildings_Draw #(parameter width_building=80)(
input					clk,
input					resetN,
input	signed [31:0]	pxl_x,
input	signed [31:0]	pxl_y,
input signed [31:0] 	topLeft_x_1,
input	signed	[31:0]	topLeft_y_1,
input signed [31:0] 	topLeft_x_2,
input	signed 	[31:0]	topLeft_y_2,

input		[31:0]	height_window,
input 				collision_building_1,
input 				collision_building_2,
output 	reg	[3:0]		Red_level,
output 	reg	[3:0]		Green_level,
output 	reg	[3:0]		Blue_level,
output 	reg				drawing_building_1,
output 	reg				drawing_building_2,
output 	reg				destructed_building_1,
output 	reg 				destructed_building_2

);

wire		in_building_1; 
wire		in_building_2; 
wire	[31:0]	offset_x_building_1;
wire	[31:0]	offset_y_building_1;
wire	[31:0]	offset_x_building_2;
wire	[31:0]	offset_y_building_2;

logic[0:79][0:79][11:0] Bitmap = {
{12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h76F,12'h76F,12'h87F,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'h98F,12'h76F,12'h75F,12'h65F,12'h65F,12'h76F,12'h76F,12'h87F,12'hA8F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h75F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'h76F,12'h66F,12'h76F,12'h76F,12'h76F,12'h66F,12'h76F,12'h76F,12'h76F,12'h75F,12'h76F,12'h77F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'h98F,12'h87F,12'h76F,12'h65F,12'h65F,12'h66F,12'h76F,12'h87F,12'h98F,12'hA9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'h98F,12'h65F,12'h65F,12'h66F,12'h76F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h75F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h76F,12'hCAF,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'hCAF,12'hB9F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h76F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hBAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hBAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h76F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hA9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hBAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hA9F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hB9F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h55F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hA8F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hBAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hA8F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h66F,12'h65F,12'h55F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h66F,12'h43F,12'hCAF,12'h43F,12'h43F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h54F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h65F,12'h66F},
{12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h87F,12'hCAF,12'h76F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h44F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h44F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h44F,12'h54F,12'h54F,12'h54F,12'h54F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'h87F,12'h98F,12'h98F,12'h98F,12'h98F,12'h98F,12'h98F,12'h98F,12'h97F,12'h87F,12'h87F,12'h87F,12'hA8F,12'hCAF,12'hCAF,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hA8F,12'h97F,12'h86F,12'h86F,12'h87F,12'h97F,12'hA8F,12'hB9F,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'hB9F,12'hA8F,12'h87F,12'h76F,12'h86F,12'h97F,12'hA8F,12'hB9F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'h97F},
{12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hBAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h98F,12'hCAF,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hA9F,12'hCAF,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hB9F,12'hCAF,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h43F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h98F,12'hCAF,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h64F,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h43F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hA8F,12'hCAF,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h53F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h43F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hA9F,12'hCAF,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h86F,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h55F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h44F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h76F,12'hCAF,12'hCAF,12'h43F,12'h66F},
{12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'h43F,12'hB9F,12'hA8F,12'h43F,12'h43F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h55F,12'h44F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'h54F,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h54F,12'h76F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h54F,12'h65F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h43F},
{12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h43F,12'h43F,12'h33F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h65F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h65F,12'h43F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hDAF,12'hCAF,12'hCAF,12'hDAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'h66F,12'h66F,12'h66F,12'h76F,12'h98F,12'hCAF,12'hCAF,12'hCAF,12'h66F,12'h66F,12'h76F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h76F,12'h75F,12'h76F,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hB9F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hA9F,12'h98F,12'h87F,12'h76F,12'h76F,12'h76F,12'h76F,12'h86F,12'h87F,12'hA9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'h87F,12'h76F,12'h66F,12'h66F,12'h66F,12'h66F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h87F,12'hCAF,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h65F,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h76F,12'hCAF,12'h97F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h54F,12'hCAF,12'h54F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h76F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h44F,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h55F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h44F,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h55F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hA8F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h55F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h44F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hA8F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h54F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h54F,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h43F,12'hCAF,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h66F,12'h65F,12'h65F,12'h65F,12'h54F,12'h43F,12'hCAF,12'h54F,12'h54F,12'h54F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h55F,12'h54F,12'h54F,12'h54F,12'h54F,12'h55F,12'hCAF,12'h43F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h43F,12'hCAF,12'h65F,12'h55F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h54F,12'h54F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h54F,12'h54F,12'h44F,12'hCAF,12'h44F,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h55F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h76F,12'hCAF,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h87F,12'hCAF,12'hB9F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h97F,12'hCAF,12'hB9F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hB9F,12'hB9F,12'hB9F,12'hC9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'h66F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h75F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'hA9F,12'hCAF,12'hCAF,12'hB9F,12'h98F,12'h87F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h86F,12'h87F,12'h98F,12'hA9F,12'hBAF,12'hCAF,12'hCAF,12'hA8F,12'h76F,12'h66F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'hCAF,12'hCAF,12'hCAF,12'h87F,12'h76F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h76F,12'h86F,12'hA8F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F},
{12'h65F,12'h65F,12'h66F,12'hCAF,12'h98F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h54F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'hCAF,12'h97F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h44F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'hCBF,12'h87F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h44F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hBAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h66F,12'hCAF,12'h87F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h66F,12'hCAF,12'h86F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h55F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h98F,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'hCBF,12'h76F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h55F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h55F,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hB9F,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h55F,12'h54F,12'h54F,12'h54F,12'hCAF,12'h65F,12'h54F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h54F,12'h54F,12'hCAF,12'h43F,12'h43F,12'h55F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h55F,12'h44F,12'h43F,12'h43F,12'hCAF,12'h54F,12'h43F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h55F,12'h44F,12'hCAF,12'h97F,12'h43F,12'h43F,12'h44F,12'h54F,12'h55F,12'h55F,12'h55F,12'h55F,12'h54F,12'h54F},
{12'h43F,12'h44F,12'h54F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h76F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h65F,12'hCAF,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h65F,12'hCAF,12'hCAF,12'h44F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h44F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'h76F,12'h65F,12'h65F,12'h65F,12'h76F,12'h76F,12'h86F,12'h87F,12'h98F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hA8F,12'h97F,12'h86F,12'h76F,12'h76F,12'h76F,12'h76F,12'h86F,12'h97F,12'hA8F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hA9F,12'hB9F,12'hB9F,12'hBAF,12'hBAF,12'hBAF,12'hBAF,12'hBAF,12'hBAF,12'hB9F,12'hB9F,12'hB9F,12'hB9F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'hB9F,12'hB9F,12'hB9F,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hB9F,12'hB9F,12'hB9F,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hA8F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hB9F,12'hCAF,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h76F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h75F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h54F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h76F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h55F,12'h66F},
{12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h54F,12'h54F,12'h54F,12'hCAF,12'h65F,12'h54F,12'h54F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h55F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h54F,12'h44F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h54F,12'h98F,12'hCAF,12'h43F,12'h55F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h54F},
{12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h65F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h65F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h54F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'h66F,12'h65F,12'h65F,12'h76F,12'h87F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hA8F,12'h97F,12'h87F,12'h76F,12'h76F,12'h76F,12'h76F,12'h76F,12'h87F,12'h87F,12'h98F,12'hA9F,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hA8F,12'h87F,12'h86F,12'h76F,12'h66F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'hCAF,12'hCAF,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h65F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h66F,12'hCAF,12'h98F,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hA8F,12'hCAF,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h97F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h98F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hBAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hA8F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'hA9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h55F,12'hB9F,12'hCAF,12'h55F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h87F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h55F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h54F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h54F,12'hCAF,12'h43F,12'h44F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h66F,12'h65F,12'h66F,12'h65F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h65F,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h55F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h66F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h55F,12'h65F,12'h65F,12'h66F},
{12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'h87F,12'h43F,12'h43F,12'h43F,12'h43F,12'h44F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hB9F,12'hB9F,12'hB9F,12'hB9F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'hB9F,12'hB9F,12'hB9F,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'h98F,12'h86F,12'h76F,12'h76F,12'h66F,12'h65F,12'h65F,12'h76F,12'h76F,12'h76F,12'h86F,12'h86F,12'h86F,12'h97F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hDAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCBF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hB9F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h54F,12'hCAF,12'h75F,12'h66F,12'h65F,12'h66F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'hCAF,12'h76F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hB9F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h44F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h97F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h98F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h54F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h76F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hA8F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h54F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h43F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hB9F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h76F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h54F,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h44F,12'h65F},
{12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h43F,12'hCAF,12'h44F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hC9F,12'hCAF,12'h43F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'hCAF,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h55F,12'h54F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h76F,12'hCAF,12'h43F,12'h55F},
{12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h44F,12'hCAF,12'h65F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h43F,12'h54F,12'h65F,12'h65F,12'h55F,12'h44F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hC9F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'h76F,12'h43F,12'h43F,12'h43F,12'h44F,12'h44F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h43F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'h87F,12'h65F,12'h64F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h65F,12'h65F,12'h65F,12'h66F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'h97F,12'h76F,12'h65F,12'h54F,12'h54F,12'h64F,12'h64F,12'h65F,12'h75F,12'h76F,12'h87F,12'hA9F,12'hCAF,12'hCAF,12'hCAF,12'hA9F,12'h65F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hB9F,12'hA9F,12'hA8F,12'hA8F,12'hA8F,12'hB9F,12'hB9F,12'hB9F,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'hB9F,12'hBAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h76F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'hCAF,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h87F,12'hCAF,12'h86F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h54F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hB9F,12'h75F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h64F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'hCAF,12'h44F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h76F,12'hCAF,12'h55F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h44F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h86F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h54F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h54F,12'hCAF,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h65F,12'h66F,12'h66F,12'h65F,12'h66F,12'h54F,12'hCAF,12'h43F,12'h55F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h66F,12'h66F,12'h66F,12'h65F,12'hA8F,12'hCAF,12'h43F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'hCAF,12'h55F,12'h54F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h65F,12'h65F,12'h44F,12'hCAF,12'h54F,12'h66F,12'h66F,12'h66F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h66F,12'h65F,12'h66F,12'h55F,12'h54F,12'hCAF,12'h54F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F,12'h65F},
{12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'hB9F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hCAF,12'h43F,12'h43F,12'h43F,12'h54F,12'h65F,12'h65F,12'h55F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'h43F,12'hCAF,12'hA9F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'hCAF,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h55F,12'hCAF,12'h55F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F,12'h54F},
{12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'h86F,12'h65F,12'h54F,12'h44F,12'h44F,12'h44F,12'h54F,12'h54F,12'h65F,12'h75F,12'h76F,12'hB9F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hA8F,12'h76F,12'h65F,12'h65F,12'h55F,12'h55F,12'h55F,12'h76F,12'h76F,12'h76F,12'h66F,12'h65F,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hCAF,12'hBAF,12'hBAF,12'hBAF}};


localparam TRANSPERENT = 12'hFFF;


assign in_building_1 = (pxl_x >= topLeft_x_1) && (pxl_x <= topLeft_x_1+width_building) &&( (pxl_y < topLeft_y_1) || (pxl_y > topLeft_y_1+height_window));
assign in_building_2 = (pxl_x >= topLeft_x_2) && (pxl_x <= topLeft_x_2+width_building) &&( (pxl_y < topLeft_y_2) || (pxl_y > topLeft_y_2+height_window));

assign offset_x_building_1 = pxl_x - topLeft_x_1;
assign offset_y_building_1 = pxl_y;
assign offset_x_building_2 = pxl_x - topLeft_x_2;
assign offset_y_building_2 = pxl_y;


always @(posedge clk or negedge resetN) begin
	if (!resetN) begin
		drawing_building_1<=0;
		drawing_building_2<=0;
		Red_level <= 4'hF;
		Green_level <= 4'hF;
		Blue_level <= 4'hF;
		destructed_building_1<=0;
		destructed_building_2<=0;
		
	end
	else begin
		drawing_building_1 <= 0;
		drawing_building_2 <= 0;
		
		if (destructed_building_1==0 && collision_building_1==1 && topLeft_x_1>-width_building) begin
			destructed_building_1<=1;
			
			
		
		end
		if (destructed_building_1==1 && topLeft_x_1<=-width_building) begin// fix to else?
			destructed_building_1<=0;
			

		end
		if (destructed_building_2==0 && collision_building_2==1 && topLeft_x_2>-width_building) begin
			destructed_building_2<=1;
			
		
		end
		if (destructed_building_2==1 && topLeft_x_2<=-width_building) begin //fix to else?
			destructed_building_2<=0;

		end
		if ((in_building_1) && (Bitmap[offset_y_building_1][offset_x_building_1]!=TRANSPERENT)&& !destructed_building_1) begin
			
			drawing_building_1 <= 1;
			Red_level <= Bitmap[{offset_y_building_1}%80][offset_x_building_1] [11:8];
			Green_level <= Bitmap[{offset_y_building_1}%80][offset_x_building_1] [7:4];
			Blue_level <= Bitmap[{offset_y_building_1}%80][offset_x_building_1] [3:0];
		end
		if ((in_building_2) && (Bitmap[offset_y_building_2][offset_x_building_2]!=TRANSPERENT) && !destructed_building_2) begin
			
			drawing_building_2 <= 1;
			Red_level <= Bitmap[{offset_y_building_2}%80][offset_x_building_2] [11:8];
			Green_level <= Bitmap[{offset_y_building_2}%80][offset_x_building_2] [7:4];
			Blue_level <= Bitmap[{offset_y_building_2}%80][offset_x_building_2] [3:0];
		end 
			
			
		
	end
end
endmodule