module light_state(
input clk,
input resetN,
input [1:0] light_num,
input [31:0] pxl_x,
input [31:0] pxl_y,
output reg draw_state_light,
output reg [31:0] red_state_light,
output reg [31:0] green_state_light,
output reg [31:0] blue_state_light,
output reg restart_light,
output reg [31:0] charging_right,
output reg [31:0] counter
);



wire [3:0] checker;


logic[0:39][0:39][11:0] Bitmap= {
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hDDD,12'hBBB,12'h888,12'h888,12'h788,12'h788,12'h778,12'h566,12'h555,12'h333,12'h000,12'hCCC},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hAAA,12'h777,12'h777,12'h777,12'h777,12'h667,12'h667,12'h556,12'h223,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h220,12'h550,12'h760,12'h660,12'h860,12'h540,12'h000,12'h000,12'hDDD,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'h777,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h100,12'h430,12'h540,12'h650,12'h660,12'h760,12'h870,12'h870,12'hBA0,12'hFD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hED0,12'h000,12'h111,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'h222,12'h000,12'h000,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFE0,12'hFF0,12'hCB0,12'h000,12'h333,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'h550,12'hFF0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFF0,12'hBA0,12'h000,12'h666,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hDDD,12'h000,12'h000,12'hCA0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFF0,12'h980,12'h000,12'hAAA,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'h888,12'h000,12'h000,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h870,12'h000,12'hCCC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'h444,12'h000,12'h220,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h650,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'h111,12'h000,12'h870,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h550,12'h112,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'h000,12'h000,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h220,12'h000,12'h779,12'h345,12'h001,12'h000,12'h000,12'h111,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hDDD,12'h000,12'h110,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hEC0,12'h000,12'h444,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'h777,12'h000,12'h660,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFF0,12'hCB0,12'h000,12'h555,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'h333,12'h000,12'hCB0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hCA0,12'h000,12'h777,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'h000,12'h000,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hCB0,12'h000,12'h999,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hEEE,12'h000,12'h660,12'hFD0,12'hB90,12'h660,12'h760,12'h650,12'h881,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hBA0,12'h000,12'hBBB,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hBBB,12'h000,12'h223,12'h668,12'h667,12'h889,12'h223,12'h000,12'hDC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hBA0,12'h000,12'hCCC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h100,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hBA0,12'h000,12'hEEE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h777,12'h000,12'h880,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hA90,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hAAA,12'h777,12'hBBB,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h000,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h980,12'h000,12'h002,12'h000,12'h000,12'h430,12'h320,12'h000,12'h000,12'h666,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDDD,12'h000,12'h650,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hED0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hBA0,12'h000,12'h000,12'hDDD,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h555,12'h000,12'hDC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFE0,12'hFF0,12'h540,12'h000,12'h111,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h110,12'hFF0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h000,12'h000,12'h666,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'h999,12'h000,12'hA90,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDC0,12'h000,12'h000,12'hCCC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'h222,12'h000,12'hFD0,12'h870,12'h650,12'h540,12'h330,12'h000,12'hDC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h870,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hCCC,12'h000,12'h444,12'h667,12'h667,12'hBCC,12'hFFF,12'hBBC,12'h000,12'hFF0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h330,12'h000,12'h666,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h233,12'h650,12'hFF0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFF0,12'hFD0,12'h000,12'h000,12'hBBB,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hFE0,12'hFE0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFE0,12'hFF0,12'h980,12'h000,12'h011,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h777,12'h210,12'hFF0,12'hFE0,12'hFE0,12'hFE0,12'hFE0,12'hFE0,12'hFE0,12'hFF0,12'h440,12'h000,12'h555,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h980,12'hFF0,12'hFE0,12'hFE0,12'hFE0,12'hFE0,12'hFF0,12'hFE0,12'h000,12'h000,12'hDDD,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'h000,12'hFE0,12'hFE0,12'hFE0,12'hFE0,12'hFE0,12'hFF0,12'hCB0,12'h000,12'h112,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h556,12'h430,12'hFF0,12'hFE0,12'hFE0,12'hFE0,12'hFF0,12'h760,12'h000,12'h777,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hCB0,12'hFE0,12'hFE0,12'hFE0,12'hFF0,12'h220,12'h000,12'hDDD,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hAAA,12'h000,12'hFF0,12'hFE0,12'hFF0,12'hED0,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h333,12'h440,12'hFF0,12'hFF0,12'hB90,12'h000,12'h666,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'hEC0,12'hFF0,12'h550,12'h000,12'hCCC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h667,12'h110,12'hFF0,12'h000,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h000,12'h550,12'h000,12'h555,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'h000,12'h000,12'hBBC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h555,12'h000,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h444,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF}};

localparam TRANSPERENT = 12'hFFF;
localparam divider_recharge = 32'd999_999_999;
assign checker[0]=(pxl_x >=500) && (pxl_x<620) &&( pxl_y<60 )&& (pxl_y>=20) && (Bitmap[pxl_y-20][{pxl_x-500}%40]!=TRANSPERENT);
assign checker[1]=(pxl_x >=540) && (pxl_x<620 )&& (pxl_y<60 )&& (pxl_y>=20)&& (Bitmap[pxl_y-20][{pxl_x-540}%40]!=TRANSPERENT);
assign checker[2]=(pxl_x >=580 )&& (pxl_x<620 )&& (pxl_y<60) && (pxl_y>=20) && (Bitmap[pxl_y-20][{pxl_x-580}%40]!=TRANSPERENT);
assign checker[3]=(pxl_x >=charging_right) && (pxl_x<620) &&( pxl_y<60 )&& (pxl_y>=20) &&( Bitmap[pxl_y-20][{pxl_x-500}%40]!=TRANSPERENT);
always @(posedge clk or negedge resetN) begin
	if (!resetN) begin
		draw_state_light<=0;
		red_state_light<=4'hF;
		green_state_light<=4'hF;
		blue_state_light<=4'hF;
		counter<=0;
		charging_right<=620;
		restart_light<=0;

		
	end
	else begin
		if (light_num==2'b11) begin
			restart_light<=0;
			
			if (checker[0]) begin
				draw_state_light<=1;
				red_state_light<=Bitmap[pxl_y-20][{pxl_x-500}%40][11:8];
				green_state_light<=Bitmap[pxl_y-20][{pxl_x-500}%40][7:4];
				blue_state_light<=Bitmap[pxl_y-20][{pxl_x-500}%40][3:0];
			end
			else begin
				draw_state_light<=0;
							
			end 
		end
		else if (light_num==2'b10) begin		
			if (checker[1]) begin
				draw_state_light<=1;
				red_state_light<=Bitmap[pxl_y-20][{pxl_x-540}%40][11:8];
				green_state_light<=Bitmap[pxl_y-20][{pxl_x-540}%40][7:4];
				blue_state_light<=Bitmap[pxl_y-20][{pxl_x-540}%40][3:0];
			end
			else begin
				draw_state_light<=0;
							
			end
		end
		else if (light_num==2'b01) begin
			if (checker[2]) begin
				draw_state_light<=1;
				red_state_light<=Bitmap[pxl_y-20][{pxl_x-580}%40][11:8];
				green_state_light<=Bitmap[pxl_y-20][{pxl_x-580}%40][7:4];
				blue_state_light<=Bitmap[pxl_y-20][{pxl_x-580}%40][3:0];

							
			end
			else begin
				draw_state_light<=0;
								
			end 
		end
		else if (light_num==0) begin
			if (charging_right>=500) begin//not yet reached end
				if (counter>divider_recharge) begin //start moving
					counter<=0;
					charging_right<=charging_right-1;
					
					if ((pxl_x >=charging_right) && (pxl_x<620) &&( pxl_y<60 )&& (pxl_y>=20) &&( Bitmap[pxl_y-20][{pxl_x-500}%40]!=TRANSPERENT)) begin
						draw_state_light<=1;
						red_state_light<=Bitmap[pxl_y-20][{pxl_x-500}%40][11:8];
						green_state_light<=Bitmap[pxl_y-20][{pxl_x-500}%40][7:4];
						blue_state_light<=Bitmap[pxl_y-20][{pxl_x-500}%40][3:0];

								
					end 
					else begin
						draw_state_light<=0;
					end
				end
				else begin
					counter<=counter+1;
				end
			end
			else begin
				restart_light=1;
				charging_right<=620;
				counter<=0;
				
			end
			
			
		end
			
		
		
		
	end
	
end
endmodule