module gameover (
input clk,
input resetN,

input [31:0] pxl_x,
input [31:0] pxl_y,
output [31:0] red_gameover,
output [31:0] green_gameover,
output [31:0] blue_gameover);

logic[0:39][0:39][11:0] GAMEOVER1={
{12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122},
{12'h111,12'h112,12'h111,12'h112,12'h112,12'h122,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h122,12'h222,12'h222,12'h222,12'h222,12'h222},
{12'h111,12'h111,12'h112,12'h122,12'h122,12'h122,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h234,12'h234,12'h233,12'h222,12'h223,12'h223,12'h223,12'h222,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h234,12'h234,12'h233,12'h222,12'h223,12'h223,12'h223,12'h223},
{12'h111,12'h112,12'h122,12'h122,12'h112,12'h245,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h367,12'h222,12'h233,12'h233,12'h233,12'h122,12'h5BD,12'h5CF,12'h5CE,12'h5CE,12'h5CF,12'h5CE,12'h233,12'h233,12'h233,12'h233,12'h223,12'h245,12'h5DF,12'h5CF,12'h48A,12'h122,12'h233,12'h233,12'h233,12'h233},
{12'h112,12'h122,12'h122,12'h112,12'h111,12'h245,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h367,12'h223,12'h233,12'h233,12'h233,12'h122,12'h5BD,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h233,12'h223,12'h233,12'h233,12'h233,12'h245,12'h5DF,12'h5CE,12'h48A,12'h122,12'h223,12'h233,12'h233,12'h233},
{12'h112,12'h122,12'h122,12'h245,12'h244,12'h356,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4BD,12'h367,12'h233,12'h233,12'h245,12'h355,12'h245,12'h4AB,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h356,12'h355,12'h255,12'h233,12'h233,12'h245,12'h5CF,12'h5CE,12'h49B,12'h245,12'h356,12'h244,12'h233,12'h233},
{12'h112,12'h122,12'h123,12'h5DF,12'h5DF,12'h4AC,12'h111,12'h122,12'h222,12'h223,12'h223,12'h223,12'h223,12'h233,12'h233,12'h233,12'h233,12'h49B,12'h5DF,12'h5DF,12'h244,12'h233,12'h233,12'h233,12'h233,12'h234,12'h5CE,12'h5DF,12'h5BD,12'h233,12'h233,12'h255,12'h5CF,12'h5CE,12'h5CE,12'h5CF,12'h5DF,12'h379,12'h233,12'h233},
{12'h122,12'h122,12'h223,12'h5CE,12'h5CE,12'h4AC,12'h122,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h233,12'h49B,12'h5CE,12'h5CF,12'h245,12'h234,12'h234,12'h234,12'h234,12'h244,12'h5CE,12'h5CE,12'h4BC,12'h233,12'h233,12'h355,12'h5CF,12'h5CE,12'h5CE,12'h5CE,12'h5CF,12'h378,12'h223,12'h222},
{12'h122,12'h122,12'h223,12'h5CE,12'h5CE,12'h4AC,12'h122,12'h233,12'h234,12'h356,12'h356,12'h356,12'h356,12'h367,12'h245,12'h234,12'h233,12'h49B,12'h5CE,12'h5CF,12'h245,12'h234,12'h244,12'h244,12'h244,12'h245,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h5BD,12'h49B,12'h4AC,12'h389,12'h356,12'h356},
{12'h122,12'h122,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h222,12'h233,12'h356,12'h5DF,12'h5CF,12'h5CF,12'h5CF,12'h5DF,12'h378,12'h234,12'h233,12'h49B,12'h5CE,12'h5CF,12'h245,12'h244,12'h244,12'h244,12'h244,12'h245,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h48A,12'h222,12'h222,12'h489,12'h5DF,12'h5DF},
{12'h122,12'h122,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h222,12'h233,12'h356,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CF,12'h378,12'h234,12'h233,12'h49B,12'h5CE,12'h5CF,12'h245,12'h234,12'h234,12'h234,12'h234,12'h244,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h49A,12'h233,12'h233,12'h48A,12'h5DF,12'h5DF},
{12'h122,12'h122,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h223,12'h233,12'h245,12'h48A,12'h489,12'h4AC,12'h5CE,12'h5CF,12'h378,12'h234,12'h234,12'h49B,12'h5CE,12'h5CE,12'h489,12'h478,12'h479,12'h479,12'h478,12'h479,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h49A,12'h233,12'h233,12'h367,12'h48A,12'h49A},
{12'h122,12'h122,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h222,12'h233,12'h233,12'h233,12'h222,12'h378,12'h5CF,12'h5CF,12'h378,12'h234,12'h234,12'h49B,12'h5CE,12'h5CE,12'h5CE,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5CE,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h244,12'h356,12'h5CF,12'h5CE,12'h49A,12'h233,12'h234,12'h233,12'h233,12'h233},
{12'h122,12'h122,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h222,12'h233,12'h233,12'h233,12'h233,12'h378,12'h5CF,12'h5CF,12'h378,12'h234,12'h234,12'h49B,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h244,12'h356,12'h5CF,12'h5CE,12'h49A,12'h233,12'h244,12'h234,12'h234,12'h234},
{12'h122,12'h122,12'h223,12'h5CE,12'h5CE,12'h4AC,12'h122,12'h233,12'h233,12'h233,12'h233,12'h378,12'h5CF,12'h5CF,12'h378,12'h233,12'h233,12'h49B,12'h5CE,12'h5CE,12'h48A,12'h489,12'h489,12'h489,12'h489,12'h48A,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h49A,12'h233,12'h234,12'h234,12'h234,12'h234},
{12'h122,12'h122,12'h123,12'h5CE,12'h5CE,12'h4AC,12'h122,12'h233,12'h233,12'h233,12'h233,12'h378,12'h5CF,12'h5CF,12'h378,12'h233,12'h233,12'h49B,12'h5CE,12'h5CF,12'h244,12'h233,12'h234,12'h234,12'h233,12'h244,12'h5CE,12'h5CE,12'h5BC,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h48A,12'h233,12'h234,12'h234,12'h234,12'h234},
{12'h112,12'h122,12'h123,12'h5DF,12'h5DF,12'h4AC,12'h111,12'h122,12'h122,12'h222,12'h122,12'h378,12'h5DF,12'h5DF,12'h378,12'h233,12'h233,12'h49B,12'h5CE,12'h5CF,12'h345,12'h234,12'h244,12'h244,12'h244,12'h244,12'h5CE,12'h5CE,12'h5BC,12'h233,12'h234,12'h355,12'h5CF,12'h5CE,12'h48A,12'h233,12'h234,12'h233,12'h233,12'h233},
{12'h112,12'h122,12'h122,12'h356,12'h256,12'h367,12'h49A,12'h49A,12'h49A,12'h49A,12'h49B,12'h379,12'h367,12'h367,12'h245,12'h233,12'h223,12'h49B,12'h5CE,12'h5CF,12'h245,12'h233,12'h234,12'h234,12'h234,12'h244,12'h5CE,12'h5CE,12'h5AC,12'h233,12'h233,12'h355,12'h5CF,12'h5CE,12'h48A,12'h223,12'h233,12'h233,12'h233,12'h233},
{12'h112,12'h112,12'h112,12'h112,12'h111,12'h244,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h389,12'h122,12'h223,12'h233,12'h233,12'h222,12'h49B,12'h5CE,12'h5DF,12'h244,12'h233,12'h234,12'h234,12'h234,12'h334,12'h5CE,12'h5CE,12'h5AC,12'h223,12'h233,12'h345,12'h5CF,12'h5CE,12'h48A,12'h222,12'h233,12'h233,12'h233,12'h233},
{12'h111,12'h112,12'h112,12'h112,12'h112,12'h245,12'h6DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h48A,12'h122,12'h223,12'h223,12'h233,12'h222,12'h4AB,12'h5DF,12'h5DF,12'h244,12'h233,12'h233,12'h233,12'h233,12'h234,12'h5CF,12'h5DF,12'h5BD,12'h222,12'h233,12'h355,12'h5DF,12'h5DF,12'h49A,12'h222,12'h233,12'h233,12'h233,12'h233},
{12'h111,12'h111,12'h112,12'h112,12'h112,12'h122,12'h234,12'h234,12'h234,12'h234,12'h244,12'h233,12'h122,12'h223,12'h223,12'h223,12'h222,12'h244,12'h245,12'h245,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h345,12'h345,12'h345,12'h233,12'h233,12'h233,12'h345,12'h345,12'h334,12'h223,12'h233,12'h233,12'h233,12'h233},
{12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h122,12'h122,12'h122,12'h222,12'h222,12'h223,12'h222,12'h222,12'h222,12'h223,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h333,12'h333,12'h333,12'h333,12'h233,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h233,12'h233,12'h233,12'h233,12'h233,12'h333,12'h333,12'h333,12'h333,12'h323,12'h223,12'h323,12'h323,12'h223,12'h223,12'h223},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h333,12'h333,12'h333,12'h333,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h223,12'h223},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h112,12'h122,12'h122,12'h122,12'h222,12'h222,12'h222,12'h222,12'h223,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323},
{12'h011,12'h011,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h112,12'h122,12'h222,12'h222,12'h222,12'h222,12'h222,12'h434,12'h534,12'h534,12'h534,12'h534,12'h534,12'h534,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323},
{12'h011,12'h011,12'h011,12'h011,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h212,12'h222,12'h222,12'h222,12'h222,12'hF8B,12'hF8B,12'hF8C,12'hF8C,12'hF8C,12'hF8B,12'hF8C,12'h534,12'h323,12'h222,12'h222,12'h323,12'h323,12'h222,12'h222,12'h222,12'h222},
{12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h212,12'h222,12'h222,12'h112,12'hE7A,12'hD7A,12'h846,12'h957,12'h856,12'hC69,12'hF8B,12'h434,12'h222,12'h856,12'h957,12'h222,12'h534,12'h957,12'h957,12'h957,12'h857},
{12'h000,12'h000,12'h000,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h212,12'h212,12'h222,12'h112,12'hF7B,12'hC69,12'h011,12'h111,12'h011,12'h856,12'hF8C,12'h434,12'h222,12'hE7A,12'hF8B,12'h122,12'h746,12'hF8C,12'hF8B,12'hF8B,12'hF8B},
{12'h001,12'h001,12'h000,12'h000,12'h000,12'h010,12'h011,12'h011,12'h011,12'h011,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h212,12'h212,12'h212,12'h112,12'hE7A,12'hE7A,12'hA57,12'hA58,12'hA57,12'hC69,12'hF8B,12'h434,12'h322,12'hE7A,12'hF7B,12'h222,12'h434,12'h846,12'h746,12'h746,12'h746},
{12'h000,12'h000,12'h000,12'h001,12'h001,12'h000,12'h000,12'h000,12'h001,12'h011,12'h001,12'h101,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h212,12'h212,12'h111,12'hE7A,12'hF8B,12'hF8C,12'hF8C,12'hF8C,12'hF8B,12'hF8C,12'h434,12'h222,12'hE7A,12'hF8B,12'h222,12'h222,12'h112,12'h112,12'h112,12'h222},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h001,12'h000,12'h000,12'h000,12'h001,12'h001,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h212,12'h111,12'hF7B,12'hD69,12'h323,12'h423,12'h433,12'h433,12'h434,12'h323,12'h322,12'hE7A,12'hF8B,12'h222,12'h645,12'hE7A,12'hD79,12'hD7A,12'hD7A},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h001,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h111,12'hF7B,12'hC69,12'h111,12'h222,12'h222,12'h222,12'h222,12'h322,12'h322,12'hE7A,12'hF8B,12'h112,12'h745,12'hF8B,12'hF7B,12'hF7B,12'hF8B},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'hF7B,12'hC69,12'h111,12'h222,12'h222,12'h222,12'h322,12'h222,12'h322,12'hE7A,12'hF8B,12'h112,12'h745,12'hF8B,12'h957,12'h222,12'h323},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h110,12'h101,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'hF7B,12'hC69,12'h111,12'h212,12'h222,12'h222,12'h322,12'h222,12'h222,12'hE7A,12'hF8B,12'h112,12'h645,12'hF8B,12'hA57,12'h433,12'h534},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h110,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'hF8B,12'hD69,12'h111,12'h212,12'h212,12'h222,12'h222,12'h222,12'h222,12'hE7A,12'hF8B,12'h111,12'h745,12'hF8B,12'hF8B,12'hF8B,12'hF8B},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h000,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'hB68,12'hA57,12'h111,12'h212,12'h212,12'h212,12'h222,12'h222,12'h222,12'hB68,12'hC69,12'h112,12'h534,12'hC69,12'hC69,12'hC69,12'hC69},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h110,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011,12'h111,12'h212,12'h212,12'h212,12'h212,12'h212,12'h212,12'h222,12'h112,12'h111,12'h222,12'h222,12'h112,12'h212,12'h212,12'h212},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h212,12'h212,12'h212,12'h212,12'h212,12'h212,12'h222,12'h222,12'h222,12'h222,12'h322,12'h322,12'h322,12'h322},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h101,12'h000,12'h111,12'h101,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111}};

logic[0:39][0:39][11:0] GAMEOVER2={
{12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h112,12'h112,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h112,12'h112,12'h112,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122},
{12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h233,12'h233,12'h233,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h122,12'h122,12'h112,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122},
{12'h223,12'h233,12'h223,12'h234,12'h234,12'h244,12'h233,12'h233,12'h233,12'h244,12'h244,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h233,12'h233,12'h233,12'h123,12'h122,12'h122,12'h122,12'h122,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h122,12'h122},
{12'h233,12'h233,12'h222,12'h5BD,12'h5CF,12'h5CF,12'h245,12'h233,12'h234,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h367,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CF,12'h49B,12'h122,12'h122},
{12'h233,12'h233,12'h222,12'h4AC,12'h5CE,12'h5CE,12'h245,12'h233,12'h244,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h367,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CF,12'h49B,12'h111,12'h222},
{12'h245,12'h356,12'h245,12'h5BD,12'h5CE,12'h5CE,12'h245,12'h233,12'h244,12'h5CE,12'h5CE,12'h5BE,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h356,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h245,12'h244,12'h245,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h49A,12'h244,12'h245},
{12'h49B,12'h5DF,12'h5CF,12'h5CE,12'h5CE,12'h5CE,12'h245,12'h234,12'h244,12'h5CE,12'h5CE,12'h5AD,12'h222,12'h233,12'h233,12'h223,12'h223,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h5CF,12'h5DF,12'h5CE,12'h111,12'h122,12'h222,12'h122,12'h122,12'h256,12'h5DF,12'h5DF},
{12'h49B,12'h5CF,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h255,12'h234,12'h245,12'h5CE,12'h5CE,12'h4BD,12'h223,12'h233,12'h233,12'h233,12'h233,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h5CE,12'h5CE,12'h5CE,12'h222,12'h223,12'h233,12'h233,12'h222,12'h356,12'h5CF,12'h5CF},
{12'h48A,12'h4AC,12'h49B,12'h5BE,12'h5CE,12'h5CE,12'h255,12'h234,12'h245,12'h5CE,12'h5CE,12'h5BD,12'h356,12'h367,12'h366,12'h356,12'h356,12'h356,12'h356,12'h356,12'h234,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h5CE,12'h5CE,12'h5CE,12'h222,12'h233,12'h233,12'h233,12'h223,12'h356,12'h5CF,12'h5CF},
{12'h367,12'h233,12'h233,12'h4AC,12'h5CE,12'h5CE,12'h355,12'h234,12'h245,12'h5CE,12'h5CE,12'h5CE,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5DF,12'h378,12'h222,12'h222,12'h122,12'h222,12'h122,12'h222,12'h122,12'h122,12'h5CE,12'h5CE,12'h5CE,12'h122,12'h233,12'h233,12'h233,12'h223,12'h356,12'h5CF,12'h5CF},
{12'h378,12'h234,12'h234,12'h4AD,12'h5CE,12'h5CE,12'h355,12'h244,12'h245,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h378,12'h222,12'h223,12'h122,12'h222,12'h222,12'h222,12'h122,12'h122,12'h5CE,12'h5CE,12'h5CE,12'h122,12'h233,12'h233,12'h233,12'h233,12'h356,12'h5CF,12'h5CF},
{12'h356,12'h234,12'h234,12'h4AD,12'h5CE,12'h5CE,12'h356,12'h244,12'h245,12'h5CE,12'h5CE,12'h5BD,12'h489,12'h48A,12'h48A,12'h48A,12'h48A,12'h489,12'h489,12'h48A,12'h255,12'h222,12'h223,12'h122,12'h222,12'h222,12'h222,12'h122,12'h222,12'h5CE,12'h5CE,12'h5CE,12'h222,12'h233,12'h233,12'h233,12'h233,12'h356,12'h5CF,12'h5CF},
{12'h234,12'h244,12'h234,12'h5AD,12'h5CE,12'h5CE,12'h255,12'h244,12'h245,12'h5CE,12'h5CE,12'h4BD,12'h223,12'h233,12'h233,12'h233,12'h233,12'h223,12'h223,12'h222,12'h222,12'h223,12'h223,12'h122,12'h222,12'h222,12'h222,12'h122,12'h222,12'h5CE,12'h5CE,12'h5CE,12'h222,12'h233,12'h233,12'h233,12'h233,12'h356,12'h5CF,12'h5CF},
{12'h234,12'h234,12'h233,12'h5AC,12'h5CE,12'h5CE,12'h355,12'h234,12'h245,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h244,12'h234,12'h234,12'h234,12'h233,12'h233,12'h233,12'h223,12'h223,12'h223,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h5CE,12'h5CE,12'h5CE,12'h222,12'h233,12'h233,12'h233,12'h233,12'h356,12'h5CF,12'h5CF},
{12'h234,12'h234,12'h233,12'h4AC,12'h5CE,12'h5CE,12'h345,12'h234,12'h245,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h244,12'h234,12'h234,12'h233,12'h233,12'h233,12'h233,12'h223,12'h223,12'h223,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h5CE,12'h5CE,12'h5CE,12'h222,12'h233,12'h233,12'h233,12'h233,12'h356,12'h5CF,12'h5CF},
{12'h234,12'h234,12'h233,12'h4AC,12'h5CE,12'h5CE,12'h345,12'h234,12'h244,12'h5CE,12'h5CE,12'h5BD,12'h233,12'h234,12'h234,12'h234,12'h233,12'h233,12'h233,12'h233,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h122,12'h5CE,12'h5CE,12'h5CE,12'h222,12'h223,12'h233,12'h233,12'h223,12'h356,12'h5CF,12'h5CF},
{12'h233,12'h234,12'h233,12'h4AC,12'h5CE,12'h5CE,12'h345,12'h233,12'h244,12'h5CE,12'h5CE,12'h5AC,12'h222,12'h233,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h5CF,12'h5DF,12'h5CF,12'h111,12'h222,12'h222,12'h222,12'h222,12'h356,12'h5DF,12'h5DF},
{12'h233,12'h233,12'h223,12'h4AC,12'h5CE,12'h5CE,12'h345,12'h233,12'h244,12'h5CE,12'h5CE,12'h5BE,12'h49A,12'h49A,12'h49A,12'h49A,12'h49A,12'h49A,12'h49A,12'h49B,12'h356,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h356,12'h356,12'h356,12'h49A,12'h49A,12'h49A,12'h49A,12'h49A,12'h489,12'h356,12'h367},
{12'h233,12'h233,12'h223,12'h5AC,12'h5CE,12'h5CE,12'h345,12'h233,12'h234,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h368,12'h122,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CF,12'h49B,12'h212,12'h222},
{12'h233,12'h233,12'h222,12'h5BD,12'h5DF,12'h5DF,12'h345,12'h233,12'h234,12'h5CF,12'h5DF,12'h5CF,12'h5CF,12'h5CF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h368,12'h212,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h4AC,12'h222,12'h223},
{12'h233,12'h233,12'h223,12'h245,12'h345,12'h345,12'h233,12'h233,12'h233,12'h345,12'h345,12'h345,12'h245,12'h245,12'h245,12'h245,12'h245,12'h244,12'h244,12'h245,12'h233,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h223,12'h222,12'h245,12'h244,12'h244,12'h244,12'h245,12'h234,12'h223,12'h223},
{12'h223,12'h233,12'h233,12'h223,12'h223,12'h223,12'h233,12'h233,12'h233,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h223},
{12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h233,12'h233,12'h233,12'h223,12'h233,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223},
{12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h323,12'h223,12'h223,12'h223,12'h223},
{12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h223},
{12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h222,12'h222,12'h222,12'h222,12'h223,12'h222,12'h223,12'h222,12'h223,12'h323,12'h322,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323},
{12'h222,12'h323,12'h323,12'h323,12'h323,12'h222,12'h222,12'h323,12'h323,12'h323,12'h222,12'h222,12'h323,12'h323,12'h323,12'h323,12'h323,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h323,12'h323,12'h323,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h323,12'h323,12'h222,12'h222,12'h222,12'h222},
{12'h957,12'h323,12'h323,12'h323,12'h323,12'h957,12'h645,12'h323,12'h323,12'h222,12'h746,12'h957,12'h222,12'h323,12'h323,12'h323,12'h222,12'h645,12'h957,12'h857,12'h857,12'h957,12'h846,12'h222,12'h323,12'h322,12'h534,12'h957,12'h957,12'h957,12'h957,12'h957,12'h957,12'h746,12'h222,12'h434,12'h957,12'h957,12'h957,12'h957},
{12'hF9C,12'h222,12'h222,12'h323,12'h434,12'hF8C,12'hA57,12'h222,12'h323,12'h222,12'hC69,12'hF8B,12'h222,12'h323,12'h323,12'h323,12'h222,12'hA58,12'hF8C,12'hF8C,12'hF8C,12'hF8C,12'hF7B,12'h111,12'h222,12'h222,12'h746,12'hF8C,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hF8C,12'hD7A,12'h222,12'h745,12'hF8C,12'hF8B,12'hF8B,12'hF8B},
{12'h745,12'hA68,12'hA57,12'h323,12'h433,12'hF8C,12'h957,12'h222,12'h323,12'h222,12'hC69,12'hF8B,12'h222,12'h323,12'h323,12'h323,12'h222,12'h534,12'h746,12'h746,12'h746,12'h746,12'h846,12'hB68,12'h957,12'h222,12'h745,12'hF8B,12'hA57,12'h746,12'h746,12'h746,12'h846,12'h745,12'h323,12'h434,12'h846,12'h746,12'h746,12'h746},
{12'h011,12'hF8B,12'hF7B,12'h323,12'h433,12'hF8C,12'h957,12'h112,12'h222,12'h111,12'hC69,12'hF8B,12'h222,12'h323,12'h323,12'h323,12'h323,12'h222,12'h112,12'h112,12'h112,12'h111,12'h323,12'hF8C,12'hD7A,12'h112,12'h745,12'hF8C,12'h645,12'h222,12'h222,12'h222,12'h222,12'h222,12'h323,12'h323,12'h212,12'h222,12'h222,12'h222},
{12'hD69,12'hF7B,12'hE7A,12'h323,12'h433,12'hF8B,12'hE7A,12'hD79,12'hD79,12'hD79,12'hE7A,12'hF7B,12'h222,12'h322,12'h323,12'h323,12'h222,12'h956,12'hD7A,12'hD79,12'hD79,12'hD79,12'hD7A,12'hF7B,12'hD79,12'h212,12'h745,12'hF8C,12'h745,12'h222,12'hB68,12'hD7A,12'hD7A,12'hB68,12'h222,12'h635,12'hE7A,12'hD79,12'hD7A,12'hD79},
{12'hF7B,12'hF7B,12'hE7A,12'h323,12'h433,12'hF8B,12'hF7B,12'hF8B,12'hF8B,12'hF7B,12'hF7B,12'hF7B,12'h222,12'h322,12'h322,12'h322,12'h222,12'hA57,12'hF8B,12'hF7B,12'hF8B,12'hF8B,12'hF7B,12'hF7B,12'hD69,12'h212,12'h745,12'hF8C,12'h745,12'h222,12'hD79,12'hF8B,12'hF8B,12'hC69,12'h222,12'h645,12'hF8B,12'hF7B,12'hF8B,12'hF8B},
{12'h212,12'hF8B,12'hE7A,12'h323,12'h322,12'h322,12'h322,12'h322,12'h222,12'h222,12'hC69,12'hF8B,12'h222,12'h322,12'h323,12'h323,12'h222,12'h957,12'hF8B,12'h635,12'h222,12'h222,12'h423,12'hF8B,12'hD69,12'h212,12'h745,12'hF8C,12'h745,12'h322,12'h323,12'h322,12'hF7B,12'hC69,12'h222,12'h645,12'hF8B,12'h957,12'h222,12'h323},
{12'h423,12'hF8B,12'hE7A,12'h323,12'h323,12'h534,12'h534,12'h534,12'h434,12'h423,12'hC69,12'hF8B,12'h222,12'h322,12'h322,12'h322,12'h222,12'h957,12'hF8B,12'h846,12'h433,12'h434,12'h634,12'hF8B,12'hD69,12'h212,12'h745,12'hF8C,12'h846,12'h534,12'h534,12'h534,12'hF7B,12'hC69,12'h212,12'h645,12'hF8B,12'hA57,12'h433,12'h534},
{12'hF8B,12'hF8B,12'hE7A,12'h323,12'h423,12'hF8C,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'h212,12'h222,12'h322,12'h322,12'h212,12'hA57,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hD7A,12'h212,12'h745,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hF8B,12'hC69,12'h212,12'h645,12'hF8B,12'hF8B,12'hF8B,12'hF8B},
{12'hC69,12'hC69,12'hB68,12'h322,12'h323,12'hC69,12'hC69,12'hC69,12'hC68,12'hC69,12'hC69,12'hC69,12'h212,12'h222,12'h322,12'h222,12'h212,12'h846,12'hC69,12'hC68,12'hC69,12'hC69,12'hC69,12'hC69,12'hA58,12'h222,12'h635,12'hC69,12'hC69,12'hC69,12'hC69,12'hC69,12'hC69,12'hA57,12'h222,12'h534,12'hC69,12'hC69,12'hC69,12'hC69},
{12'h212,12'h212,12'h212,12'h322,12'h222,12'h212,12'h212,12'h112,12'h112,12'h112,12'h112,12'h212,12'h222,12'h222,12'h222,12'h222,12'h322,12'h212,12'h112,12'h112,12'h212,12'h212,12'h212,12'h212,12'h222,12'h322,12'h222,12'h212,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h323,12'h222,12'h222,12'h212,12'h212,12'h212},
{12'h322,12'h322,12'h322,12'h322,12'h322,12'h322,12'h322,12'h322,12'h322,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h322,12'h322,12'h322,12'h322,12'h322,12'h322,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323,12'h323},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111}};
logic[0:39][0:39][11:0] GAMEOVER3={
{12'h122,12'h122,12'h122,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h122,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122},
{12'h122,12'h122,12'h122,12'h122,12'h112,12'h112,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h223,12'h223,12'h222,12'h223,12'h223,12'h223,12'h223,12'h233,12'h223,12'h223,12'h233,12'h233,12'h223,12'h233,12'h233,12'h233,12'h223,12'h223,12'h222,12'h222,12'h222},
{12'h122,12'h122,12'h122,12'h133,12'h233,12'h233,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h233,12'h234,12'h233,12'h223,12'h223,12'h233,12'h244,12'h234,12'h234,12'h244,12'h244,12'h244,12'h244,12'h244,12'h244,12'h244,12'h244,12'h233,12'h233,12'h233,12'h234,12'h234,12'h234,12'h234,12'h234},
{12'h122,12'h122,12'h111,12'h49A,12'h5CF,12'h5DF,12'h256,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h233,12'h5CF,12'h5CF,12'h4AC,12'h122,12'h223,12'h255,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h245,12'h233,12'h222,12'h5BD,12'h5CF,12'h5CE,12'h5CE,12'h5CE},
{12'h222,12'h223,12'h112,12'h49A,12'h5CE,12'h5CF,12'h256,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h222,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h222,12'h223,12'h355,12'h5DF,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h255,12'h233,12'h223,12'h5BD,12'h5CE,12'h5CE,12'h5CE,12'h5CE},
{12'h234,12'h222,12'h122,12'h49A,12'h5CE,12'h5CF,12'h256,12'h122,12'h222,12'h222,12'h222,12'h222,12'h223,12'h222,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h223,12'h233,12'h255,12'h5CF,12'h5CE,12'h5BD,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h4AC,12'h5BD,12'h245,12'h233,12'h233,12'h5BD,12'h5CE,12'h5CE,12'h4AC,12'h4AC},
{12'h489,12'h122,12'h122,12'h49A,12'h5CE,12'h5CF,12'h356,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h223,12'h233,12'h255,12'h5CF,12'h5CE,12'h48A,12'h223,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h234,12'h233,12'h5BD,12'h5CE,12'h5BE,12'h233,12'h223},
{12'h389,12'h222,12'h122,12'h49A,12'h5CE,12'h5CF,12'h356,12'h222,12'h223,12'h223,12'h233,12'h233,12'h233,12'h233,12'h233,12'h5CE,12'h5CE,12'h4AC,12'h233,12'h233,12'h356,12'h5CF,12'h5CE,12'h48A,12'h233,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h233,12'h5BD,12'h5CE,12'h5BE,12'h234,12'h233},
{12'h389,12'h223,12'h222,12'h49A,12'h5CE,12'h5CF,12'h356,12'h222,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h5CE,12'h5CE,12'h4AC,12'h233,12'h233,12'h356,12'h5CF,12'h5CE,12'h49B,12'h356,12'h367,12'h367,12'h367,12'h367,12'h367,12'h367,12'h367,12'h245,12'h244,12'h233,12'h5BD,12'h5CE,12'h5BE,12'h367,12'h356},
{12'h489,12'h223,12'h222,12'h49A,12'h5CE,12'h5CF,12'h356,12'h222,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h5CE,12'h5CE,12'h4AC,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h5CE,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5CF,12'h5DF,12'h356,12'h234,12'h233,12'h5BD,12'h5CE,12'h5CE,12'h5CF,12'h5CF},
{12'h489,12'h223,12'h222,12'h49A,12'h5CE,12'h5CF,12'h356,12'h222,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h5CE,12'h5CE,12'h4AC,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h356,12'h234,12'h233,12'h5BD,12'h5CE,12'h5CE,12'h5CE,12'h5CE},
{12'h489,12'h223,12'h222,12'h49A,12'h5CE,12'h5CF,12'h356,12'h223,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h5CE,12'h5CE,12'h4AC,12'h233,12'h234,12'h356,12'h5CF,12'h5CE,12'h4AC,12'h48A,12'h48A,12'h48A,12'h48A,12'h48A,12'h48A,12'h48A,12'h49A,12'h245,12'h234,12'h233,12'h5BD,12'h5CE,12'h5CE,12'h48A,12'h48A},
{12'h489,12'h223,12'h222,12'h49A,12'h5CE,12'h5CF,12'h356,12'h223,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h234,12'h5CE,12'h5CE,12'h4AC,12'h233,12'h233,12'h356,12'h5CF,12'h5CE,12'h48A,12'h233,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h244,12'h244,12'h233,12'h5BD,12'h5CE,12'h5BE,12'h233,12'h233},
{12'h489,12'h223,12'h222,12'h49B,12'h5DF,12'h5DF,12'h356,12'h122,12'h222,12'h233,12'h233,12'h233,12'h223,12'h223,12'h233,12'h5CF,12'h5CF,12'h4AC,12'h233,12'h233,12'h356,12'h5CF,12'h5CE,12'h48A,12'h234,12'h244,12'h244,12'h244,12'h244,12'h244,12'h244,12'h244,12'h244,12'h234,12'h233,12'h5BD,12'h5CE,12'h5BE,12'h244,12'h233},
{12'h489,12'h223,12'h223,12'h367,12'h389,12'h379,12'h378,12'h378,12'h479,12'h233,12'h233,12'h223,12'h479,12'h378,12'h378,12'h389,12'h489,12'h378,12'h233,12'h233,12'h356,12'h5CF,12'h5CE,12'h48A,12'h234,12'h244,12'h244,12'h244,12'h244,12'h244,12'h244,12'h234,12'h234,12'h234,12'h233,12'h5BD,12'h5CE,12'h5BE,12'h234,12'h233},
{12'h389,12'h223,12'h233,12'h223,12'h222,12'h111,12'h49B,12'h5DF,12'h5DF,12'h234,12'h223,12'h122,12'h5DF,12'h5CF,12'h5CE,12'h222,12'h223,12'h233,12'h234,12'h233,12'h356,12'h5CF,12'h5CE,12'h48A,12'h233,12'h244,12'h234,12'h244,12'h234,12'h234,12'h234,12'h234,12'h234,12'h234,12'h233,12'h5BD,12'h5CE,12'h5BE,12'h234,12'h233},
{12'h489,12'h222,12'h233,12'h233,12'h233,12'h222,12'h4AB,12'h5DF,12'h5DF,12'h233,12'h222,12'h111,12'h5DF,12'h5DF,12'h5CE,12'h233,12'h233,12'h233,12'h234,12'h233,12'h356,12'h5CF,12'h5CE,12'h48A,12'h222,12'h233,12'h233,12'h233,12'h233,12'h233,12'h233,12'h223,12'h233,12'h233,12'h223,12'h5BD,12'h5CE,12'h5BE,12'h234,12'h233},
{12'h245,12'h223,12'h233,12'h233,12'h223,12'h222,12'h255,12'h367,12'h356,12'h48A,12'h49A,12'h49B,12'h356,12'h367,12'h366,12'h233,12'h233,12'h233,12'h233,12'h233,12'h355,12'h5CF,12'h5CE,12'h5BD,12'h49A,12'h49B,12'h49A,12'h49A,12'h49A,12'h49A,12'h49A,12'h49B,12'h244,12'h233,12'h222,12'h5BD,12'h5CE,12'h5BE,12'h233,12'h223},
{12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h111,12'h5BE,12'h5CF,12'h5DF,12'h212,12'h222,12'h222,12'h233,12'h233,12'h233,12'h233,12'h233,12'h355,12'h5CF,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5CE,12'h5DF,12'h245,12'h223,12'h122,12'h5BD,12'h5CE,12'h5BE,12'h233,12'h222},
{12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h111,12'h5CE,12'h5DF,12'h6EF,12'h222,12'h223,12'h223,12'h223,12'h233,12'h233,12'h233,12'h223,12'h355,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h5DF,12'h245,12'h222,12'h122,12'h5CE,12'h5DF,12'h5CF,12'h233,12'h122},
{12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h244,12'h244,12'h245,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h233,12'h245,12'h245,12'h245,12'h245,12'h245,12'h245,12'h245,12'h245,12'h245,12'h244,12'h245,12'h223,12'h222,12'h122,12'h244,12'h244,12'h234,12'h122,12'h122},
{12'h223,12'h223,12'h223,12'h223,12'h222,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h112,12'h112,12'h122,12'h122},
{12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h112,12'h112},
{12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h223,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h112,12'h112,12'h112,12'h111},
{12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h112,12'h112,12'h112,12'h112,12'h111,12'h111,12'h111,12'h111},
{12'h323,12'h323,12'h323,12'h322,12'h223,12'h223,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h433,12'h434,12'h434,12'h434,12'h434,12'h433,12'h222,12'h222,12'h222,12'h122,12'h122,12'h122,12'h112,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111},
{12'h222,12'h323,12'h323,12'h323,12'h222,12'h222,12'h222,12'h323,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h222,12'h011,12'hD79,12'hF8C,12'hF8C,12'hF8C,12'hF8C,12'hD69,12'h011,12'h112,12'h212,12'h112,12'h112,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111},
{12'h957,12'h323,12'h323,12'h222,12'h534,12'h957,12'h645,12'h222,12'h645,12'h957,12'h323,12'h222,12'h222,12'h323,12'h957,12'h635,12'h122,12'h534,12'h957,12'h956,12'h856,12'h846,12'h846,12'h846,12'h846,12'h856,12'h434,12'h111,12'h112,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111},
{12'hF8C,12'h323,12'h222,12'h222,12'h746,12'hF9D,12'hB68,12'h111,12'hB68,12'hF8C,12'h423,12'h112,12'h222,12'h434,12'hF8C,12'hA57,12'h111,12'hA57,12'hF9D,12'h534,12'h111,12'h112,12'h111,12'h000,12'h433,12'hF9D,12'h846,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011,12'h011,12'h011},
{12'h745,12'hA58,12'hA57,12'h323,12'h434,12'h846,12'h534,12'h212,12'hA58,12'hF8B,12'hB68,12'hB68,12'h222,12'h434,12'hF8B,12'h957,12'h111,12'h534,12'h846,12'h323,12'h222,12'h222,12'h212,12'hB68,12'h957,12'h745,12'h323,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011,12'h011,12'h011,12'h011},
{12'h011,12'hE7A,12'hF7B,12'h323,12'h222,12'h112,12'h222,12'h222,12'hA58,12'hF8B,12'hF8B,12'hF8C,12'h011,12'h323,12'hF8B,12'h957,12'h112,12'h212,12'h212,12'h212,12'h212,12'h111,12'h111,12'hF9D,12'hC69,12'h011,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011,12'h001,12'h001,12'h001,12'h010},
{12'hD69,12'hF7B,12'hE7A,12'h222,12'h645,12'hE7A,12'h957,12'h112,12'hA58,12'hF8B,12'h634,12'h323,12'hD7A,12'hD7A,12'hF8B,12'h957,12'h112,12'h222,12'h222,12'h212,12'h222,12'hC69,12'hD7A,12'h222,12'h322,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h101,12'h101,12'h101,12'h000,12'h000,12'h000},
{12'hF7B,12'hF7B,12'hE7A,12'h222,12'h745,12'hF8C,12'hA57,12'h111,12'hA58,12'hF8B,12'h423,12'h111,12'hF8B,12'hF8B,12'hF8B,12'h957,12'h111,12'h212,12'h212,12'h212,12'h212,12'hE7A,12'hF8B,12'h000,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h001,12'h101,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h212,12'hE7A,12'hE7A,12'h322,12'h645,12'hF8B,12'hA57,12'h111,12'hA58,12'hF8B,12'h433,12'h222,12'h222,12'h433,12'hF8B,12'h957,12'h111,12'h212,12'h212,12'h212,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h110,12'h110,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h423,12'hE7A,12'hE7A,12'h222,12'h645,12'hF8B,12'hA57,12'h111,12'hA58,12'hF8B,12'h423,12'h222,12'h212,12'h423,12'hF8B,12'h957,12'h111,12'h212,12'h212,12'h212,12'h112,12'h323,12'h423,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011,12'h110,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'hF8B,12'hF8B,12'hE7A,12'h222,12'h745,12'hF8C,12'hA57,12'h111,12'hA68,12'hF8B,12'h423,12'h212,12'h212,12'h423,12'hF8B,12'h957,12'h111,12'h212,12'h212,12'h112,12'h212,12'hF8B,12'hF8C,12'h000,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h001,12'h110,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'hC69,12'hC69,12'hB68,12'h222,12'h634,12'hD79,12'h846,12'h111,12'h846,12'hC69,12'h423,12'h222,12'h212,12'h323,12'hC69,12'h746,12'h111,12'h212,12'h212,12'h111,12'h111,12'hB68,12'hC69,12'h000,12'h111,12'h111,12'h111,12'h111,12'h111,12'h101,12'h110,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h212,12'h212,12'h212,12'h322,12'h222,12'h112,12'h212,12'h322,12'h212,12'h111,12'h212,12'h212,12'h212,12'h212,12'h111,12'h111,12'h212,12'h212,12'h111,12'h111,12'h111,12'h001,12'h000,12'h111,12'h111,12'h111,12'h111,12'h111,12'h101,12'h011,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h322,12'h322,12'h322,12'h322,12'h322,12'h322,12'h222,12'h222,12'h222,12'h222,12'h212,12'h212,12'h212,12'h212,12'h212,12'h212,12'h212,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h110,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h101,12'h111,12'h100,12'h101,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000}};
logic[0:39][0:9][11:0] GAMEOVER4={
{12'h122,12'h122,12'h122,12'h122,12'h122,12'h112,12'h111,12'h111,12'h111,12'h011},
{12'h122,12'h122,12'h122,12'h122,12'h122,12'h122,12'h112,12'h112,12'h112,12'h011},
{12'h234,12'h233,12'h233,12'h233,12'h122,12'h122,12'h122,12'h112,12'h112,12'h111},
{12'h5CE,12'h5CE,12'h5CF,12'h4BD,12'h111,12'h122,12'h122,12'h122,12'h122,12'h111},
{12'h5CE,12'h5CE,12'h5CF,12'h4BD,12'h111,12'h122,12'h122,12'h122,12'h122,12'h111},
{12'h4AC,12'h4AC,12'h4AC,12'h49B,12'h244,12'h245,12'h234,12'h112,12'h122,12'h111},
{12'h223,12'h223,12'h122,12'h234,12'h5DF,12'h5DF,12'h49B,12'h111,12'h122,12'h111},
{12'h233,12'h233,12'h222,12'h244,12'h5DF,12'h5CF,12'h49A,12'h111,12'h122,12'h111},
{12'h356,12'h356,12'h356,12'h367,12'h4AC,12'h4AB,12'h378,12'h122,12'h122,12'h111},
{12'h5CF,12'h5CF,12'h5DF,12'h5BD,12'h111,12'h122,12'h122,12'h122,12'h122,12'h111},
{12'h5CE,12'h5CE,12'h5CF,12'h5BD,12'h111,12'h222,12'h122,12'h122,12'h122,12'h111},
{12'h48A,12'h489,12'h489,12'h389,12'h377,12'h378,12'h356,12'h122,12'h122,12'h111},
{12'h233,12'h223,12'h222,12'h244,12'h5DF,12'h5DF,12'h49B,12'h111,12'h122,12'h111},
{12'h233,12'h233,12'h233,12'h244,12'h5DF,12'h5CE,12'h49A,12'h111,12'h122,12'h111},
{12'h233,12'h233,12'h223,12'h244,12'h5DF,12'h5CE,12'h48A,12'h111,12'h122,12'h111},
{12'h233,12'h233,12'h223,12'h244,12'h5DF,12'h5CE,12'h48A,12'h111,12'h122,12'h111},
{12'h233,12'h223,12'h222,12'h234,12'h5DF,12'h5CE,12'h48A,12'h111,12'h122,12'h111},
{12'h223,12'h223,12'h122,12'h234,12'h5DF,12'h5CE,12'h48A,12'h111,12'h122,12'h111},
{12'h222,12'h122,12'h122,12'h234,12'h5DF,12'h5CE,12'h48A,12'h111,12'h122,12'h111},
{12'h122,12'h122,12'h122,12'h234,12'h6EF,12'h5DF,12'h49B,12'h111,12'h112,12'h111},
{12'h122,12'h122,12'h122,12'h122,12'h234,12'h134,12'h123,12'h111,12'h111,12'h011},
{12'h122,12'h112,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011},
{12'h112,12'h112,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011},
{12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h111,12'h011,12'h011,12'h001},
{12'h111,12'h111,12'h111,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h000},
{12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h000},
{12'h011,12'h011,12'h011,12'h011,12'h011,12'h011,12'h010,12'h000,12'h000,12'h000},
{12'h011,12'h011,12'h010,12'h000,12'h000,12'h000,12'h000,12'h001,12'h001,12'h000},
{12'h000,12'h000,12'h000,12'h001,12'h001,12'h001,12'h001,12'h000,12'h000,12'h000},
{12'h001,12'h001,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000}};

always @(posedge clk or negedge resetN) begin
			if (!resetN) begin
			end 
			else begin
				if ((pxl_y >=220) && (pxl_y<260)) begin
					if ((pxl_x>=255) && (pxl_x<295)) begin
						red_gameover<= GAMEOVER1[pxl_y-220][pxl_x-255][11:8];
						green_gameover<= GAMEOVER1[pxl_y-220][pxl_x-255][7:4];
						blue_gameover<= GAMEOVER1[pxl_y-220][pxl_x-255][3:0];
					end
					else if ((pxl_x>=295) && (pxl_x<335)) begin
						red_gameover<= GAMEOVER2[pxl_y-220][pxl_x-295][11:8];
						green_gameover<= GAMEOVER2[pxl_y-220][pxl_x-295][7:4];
						blue_gameover<= GAMEOVER2[pxl_y-220][pxl_x-295][3:0];
					end
					else if ((pxl_x>=335) && (pxl_x<375)) begin
						red_gameover<= GAMEOVER3[pxl_y-220][pxl_x-335][11:8];
						green_gameover<= GAMEOVER3[pxl_y-220][pxl_x-335][7:4];
						blue_gameover<= GAMEOVER3[pxl_y-220][pxl_x-335][3:0];
					end
					else if ((pxl_x>=375) && (pxl_x<385)) begin
						red_gameover<= GAMEOVER4[pxl_y-220][pxl_x-375][11:8];
						green_gameover<= GAMEOVER4[pxl_y-220][pxl_x-375][7:4];
						blue_gameover<= GAMEOVER4[pxl_y-220][pxl_x-375][3:0];
					end
					else begin
						red_gameover<=4'h0;
						green_gameover<= 4'h0;
						blue_gameover<=4'h0;
					end
					
					
				end
				else begin
					red_gameover<=4'h0;
					green_gameover<= 4'h0;
					blue_gameover<=4'h0;
				end
			end
			
			
end
endmodule