module Bird_Draw #( height_bird=56,  width_bird=100)(
input					clk,
input					resetN,
input		[31:0]	pxl_x,
input		[31:0]	pxl_y,
input		integer 	topLeft_x_bird,
input		integer	topLeft_y_bird,


output reg	[3:0]		Red_level,
output reg	[3:0]		Green_level,
output reg	[3:0]		Blue_level,
output reg				drawing_bird);

wire	in_rectangle; 
wire	[31:0]	offset_x;
wire	[31:0]	offset_y;

logic[0:(height_bird-1)][0:(width_bird-1)][11:0] Bitmap = {
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hDDE,12'hCCE,12'hCCE,12'h99E,12'h00E,12'h11E,12'h33E,12'h66E,12'h889,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hBBD,12'hBBF,12'hBBF,12'hDDF,12'h88F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h009,12'h005,12'h88A,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEDD,12'hD99,12'hD44,12'hD55,12'hD77,12'hBCE,12'hBBF,12'hCCF,12'hCCF,12'h88F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h005,12'h007,12'h006,12'hEEE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDBC,12'hEAB,12'hF55,12'hE00,12'hE11,12'hF00,12'hB7A,12'hCCF,12'hCCF,12'hCCF,12'hDDF,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h007,12'h005,12'h003,12'h888,12'hFFE,12'hEEE,12'hEEE,12'hFEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEAA,12'hFBB,12'hF67,12'hE01,12'hE12,12'hF11,12'hC57,12'hCDF,12'hCCF,12'hCCF,12'hCCF,12'h99F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h8D9,12'hBFA,12'h7F7,12'h0F0,12'h0E0,12'h5E5,12'hDED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDAA,12'hFAB,12'hFBC,12'hE23,12'hE12,12'hF12,12'hC01,12'h89F,12'hCCF,12'hCCF,12'hCCF,12'hDDF,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'hCFA,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h3D3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDCC,12'hFAA,12'hFBB,12'hFBC,12'hE12,12'hE12,12'hF11,12'h30A,12'h12F,12'hEEF,12'hDDF,12'hBBF,12'h11F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h169,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hEEE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hE9A,12'hFBB,12'hFBB,12'hFBB,12'hE01,12'hF12,12'hE11,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hFEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDCD,12'hFBB,12'hFBB,12'hFCC,12'hF55,12'hE11,12'hF11,12'h706,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h076,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h3D3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD55,12'hF67,12'hF77,12'hF44,12'hE01,12'hE12,12'hF11,12'h20B,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00D,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hDED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hE00,12'hE11,12'hE11,12'hE11,12'hE12,12'hE12,12'hF10,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h5D5,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDBB,12'hE01,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hE11,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h0A3,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0E0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD88,12'hE01,12'hE12,12'hE12,12'hE12,12'hE12,12'hF12,12'hC12,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h076,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hFEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD67,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hF12,12'hC12,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h049,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hFEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD55,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hF12,12'hC12,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00D,12'h006,12'h00F,12'h00F,12'h00F,12'h03A,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hEEE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD55,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hF12,12'hD11,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h000,12'h000,12'h005,12'h00F,12'h02D,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hFEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD66,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h007,12'h000,12'h000,12'h000,12'h003,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hEE8,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD77,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF10,12'h00F,12'h00F,12'h00F,12'h009,12'h00C,12'h00E,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h000,12'h000,12'h870,12'hBB0,12'h860,12'h4A0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0F0,12'h0D0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hDD7,12'hEE1,12'hFF0,12'hFF0,12'hEEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD99,12'hE01,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'h20B,12'h00F,12'h00F,12'h002,12'h000,12'h000,12'h000,12'h000,12'h003,12'h008,12'h00C,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00C,12'h330,12'hFE0,12'hFD0,12'hFF0,12'hFF0,12'hFF0,12'h5D0,12'h0F0,12'h0F0,12'h0F0,12'h4E4,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEED,12'hDD7,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEDD,12'hE00,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'h608,12'h00F,12'h00F,12'h00F,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h110,12'h550,12'h662,12'h667,12'h11C,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h436,12'hFD0,12'hEC0,12'hEC0,12'hED0,12'hFF0,12'hFF0,12'hDE0,12'h1E0,12'h0F0,12'h8E8,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hEE7,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD01,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'hB13,12'h00F,12'h00F,12'h00F,12'h00F,12'h000,12'h000,12'h000,12'h000,12'hDD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h994,12'h22B,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'hB92,12'hFD0,12'hEC0,12'hEC0,12'hEC0,12'hFD0,12'hFF0,12'hFF0,12'h7D0,12'hDDF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEA,12'hEE2,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD44,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF10,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h000,12'h000,12'h430,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h994,12'h11C,12'h00F,12'h00F,12'h00F,12'hDA0,12'hFC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFE0,12'hEED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hDD7,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDBB,12'hE01,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'h806,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h000,12'h100,12'hFD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'h667,12'h00F,12'h0C0,12'hDC0,12'hFC0,12'hEC0,12'hEC0,12'hEC0,12'hEB0,12'hFF0,12'hFF0,12'hFF0,12'hDD8,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hDD4,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD01,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF10,12'h00E,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h002,12'hCA0,12'hEC0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hAE0,12'h0D0,12'hBB0,12'hFC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hEE5,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hDD4,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE1,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD99,12'hE01,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'hC13,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h226,12'hFE0,12'hEC0,12'hED0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hBD0,12'hCB0,12'hDB0,12'hDB0,12'hDC0,12'hED0,12'hDD0,12'hDD0,12'hDD0,12'hEE0,12'hDD2,12'hEE6,12'hDDB,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hDD6,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE2,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hD22,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'h806,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h22B,12'hFD0,12'hFC0,12'hEC0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hDD5,12'hEEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hDDA,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE2,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hE00,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'h815,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'hCA1,12'hFD0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hEE6,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE2,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hDDC,12'hEEA,12'hEE7,12'hDD5,12'hDD8,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hECC,12'hE00,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hE12,12'hF11,12'hC12,12'h00D,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h00F,12'h548,12'hFD0,12'hFC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD6,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hEE2,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFD0,12'hEC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hEE2,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hDD9,12'hEE4,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDCC,12'hE00,12'hE11,12'hE12,12'hE12,12'hE12,12'hE12,12'hE02,12'hE02,12'hE10,12'hA33,12'h448,12'h666,12'h885,12'h995,12'h556,12'h33A,12'h33A,12'hBA0,12'hEC0,12'hEC0,12'hEC0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD7,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hEE8,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hED0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFE0,12'hFF0,12'hEE2,12'hFFF,12'hEEC,12'hEE6,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEEC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hD23,12'hE00,12'hF02,12'hE02,12'hD51,12'hDB0,12'hEF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hCA0,12'hDB0,12'hEC0,12'hEC0,12'hFD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEED,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hEEE,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hED0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDAC,12'hD60,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hEB0,12'hCA0,12'hEB0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE1,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hEE1,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEEB,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hEF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFD0,12'hDB0,12'hCA0,12'hEB0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hEEC,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hDD9,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFE0,12'hFD0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDDA,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEB,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD0,12'hEE0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFD0,12'hDB0,12'hCA0,12'hDB0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD0,12'hFFF,12'h883,12'hFF0,12'hFF0,12'hEE5,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hCB1,12'hEC0,12'hEC0,12'hEC0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFD0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hEE0,12'hEE1,12'hCA3,12'hB88,12'hC98,12'hCA9,12'hCBA,12'hDCC,12'hDDA,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h550,12'h001,12'h110,12'hFF0,12'hFF0,12'hEE0,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hDD6,12'hFF0,12'hFF0,12'hED0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB0,12'hDDA,12'hEFF,12'hEB0,12'hEC0,12'hEC0,12'hFD0,12'hFF0,12'hED0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEC1,12'hB75,12'hB74,12'hA64,12'hA63,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h220,12'h000,12'h110,12'hFF0,12'hFF0,12'hFF0,12'hEEE,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hEEF,12'hEE0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB3,12'hFFF,12'hFFF,12'hFFF,12'hDB0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFE0,12'hFF0,12'hFF0,12'hFD0,12'hED0,12'hEC0,12'hEC0,12'hB81,12'h962,12'h853,12'h853,12'h733,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h110,12'h000,12'h220,12'hFF0,12'hFF0,12'hFF0,12'hDDB,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hDB5,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEB0,12'hDC9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDB2,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB0,12'hDC7,12'hCB4,12'hEC0,12'hEC0,12'hEC0,12'hFD0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hFC0,12'hEC0,12'h742,12'h733,12'hBB0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h330,12'h000,12'h660,12'hFF0,12'hFF0,12'hFF0,12'hEE9,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hEB0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB0,12'hEED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDC6,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEB0,12'hDB4,12'hDDC,12'hFFF,12'hFFF,12'hEDA,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB0,12'hDC4,12'hCBA,12'hEEE,12'hEEC,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hDD0,12'hDD0,12'hDD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEB0,12'hE10,12'hE00,12'hE00,12'hD70,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h880,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE2,12'hEEC,12'hEEF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDC5,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB1,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEDD,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB0,12'hDC5,12'hEEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDDD,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB0,12'hDC5,12'hEDC,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD0,12'hEE0,12'hFF0,12'hEE0,12'hEE0,12'hEE0,12'hDD0,12'hEE0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hE80,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hE10,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'h993},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hDB0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDB0,12'hEC0,12'hEB0,12'hDB4,12'hEEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDB0,12'hEC0,12'hEC0,12'hDB0,12'hDC8,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD8,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD0,12'hFF0,12'hEE0,12'hDD0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hEE0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEF0,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hE80,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE4},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDC7,12'hEC0,12'hEC0,12'hEC0,12'hDC5,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDC8,12'hDB0,12'hEED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDB3,12'hDB0,12'hDDA,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hCC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hD90,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hD20,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE6},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDB0,12'hEC0,12'hDC7,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD8,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hCC0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hE80,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hE10,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEEB},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD9,12'hDC6,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hDD0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hED0,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hE60,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDC1,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD9,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hEE0,12'hDD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hD40,12'hF00,12'hF00,12'hF00,12'hF00,12'hF00,12'hE00,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hD95,12'hD78,12'hEEA,12'hDD6,12'hDD6,12'hEEC,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEE1,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hDD0,12'hFF0,12'hDD0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hD60,12'hF00,12'hF00,12'hF00,12'hE10,12'hEF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hD76,12'hDBD,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD5,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hEE0,12'hFF0,12'hEE0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDC0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD6,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDD0,12'hEE0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hDD0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEEE,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE1,12'hEEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD3,12'hFF0,12'hFF0,12'hFF0,12'hED0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hDB0,12'hFD0,12'hEE0,12'hFF0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hDD9,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEF,12'hFF0,12'hFF0,12'hFF0,12'hEC0,12'hDB3,12'hEEA,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hDB0,12'hEC0,12'hEC0,12'hEC0,12'hDC0,12'hFF0,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE3,12'hDDA,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEE8,12'hFF0,12'hFF0,12'hEC0,12'hEB0,12'hEED,12'hFFF,12'hEEF,12'hDD5,12'hEE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hDC0,12'hCA0,12'hCA0,12'hDB0,12'hCB0,12'hDB0,12'hB90,12'hDB0,12'hDB0,12'hFE0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hFF0,12'hEE0,12'hDD2,12'hEE7,12'hDDB,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEE2,12'hFF0,12'hFF0,12'hEC0,12'hDB5,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEB,12'hDD6,12'hEE3,12'hEE1,12'hDD0,12'hEE2,12'hDD1,12'hDC0,12'hDB0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB1,12'hFFF,12'hFFF,12'hEEF,12'hDDD,12'hEDC,12'hEEB,12'hEE9,12'hDD8,12'hDD7,12'hDD7,12'hDD5,12'hDD5,12'hDD5,12'hDD5,12'hDD7,12'hDD7,12'hEE9,12'hEEA,12'hEEB,12'hEED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDD0,12'hFF0,12'hEC0,12'hDB0,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDB5,12'hEB0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hEC0,12'hDB3,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hDE0,12'hEF0,12'hDB0,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEEE,12'hDC8,12'hDC4,12'hDC4,12'hDC6,12'hEED,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDDC,12'hFF0,12'hCC0,12'hFEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF},
{12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEED,12'hEE7,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF}};
localparam TRANSPERENT = 12'hFFF;
	

assign in_rectangle = (pxl_x >= topLeft_x_bird) && (pxl_x < topLeft_x_bird+width_bird) && (pxl_y >= topLeft_y_bird) && (pxl_y < topLeft_y_bird+height_bird);
assign offset_x = pxl_x - topLeft_x_bird;
assign offset_y = pxl_y - topLeft_y_bird;
always @(posedge clk or negedge resetN) begin
	if (!resetN) begin
		drawing_bird<=0;
		Red_level <= 4'hF;
		Green_level <= 4'hF;
		Blue_level <= 4'hF;
	end
	else begin
		drawing_bird <= 0;
		if ((in_rectangle) && (Bitmap[offset_y][offset_x]!=TRANSPERENT)) begin
			
			drawing_bird <= 1;
			Red_level <= Bitmap[offset_y][offset_x] [11:8];
			Green_level <= Bitmap[offset_y][offset_x] [7:4];
			Blue_level <= Bitmap[offset_y][offset_x] [3:0];
		end
			
			
		
	end
end


endmodule