module Background_Draw #(parameter screen_size=640)(
input [31:0] pxl_x,
input [31:0] pxl_y,
input clk, 
output background_drawing, 
output reg [3:0] Blue_background,
output reg [3:0] Green_background,
output reg [3:0] Red_background);


logic[0:79][0:79][11:0] Bitmap={
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h6EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h6EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h8EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7DF,12'hFFF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h8EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h8EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'h7EF,12'hCEF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7CF,12'hFFF,12'hFFF,12'h7EF,12'hBEF,12'h7DF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7FF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h8EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h8EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h7EF,12'h7FF,12'h7EF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'h7EF,12'h7EF,12'h7EF,12'h8EF,12'hFFF,12'hFFF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'h7FF,12'h7EF,12'h7EF,12'hEFF,12'hFFF,12'hEFF,12'h7EF,12'h7EF,12'hEFF,12'hFFF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7FF,12'h8DF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'h9DF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h7EF,12'h8EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'h8EF,12'h7EF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'h8EF,12'h8EF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'h7EF,12'hFFF,12'hFFF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hEFF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h7DF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'h9DF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h8FF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'h7EF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hEEF,12'hFFF,12'h7FF,12'h7EF,12'h7EF,12'h7EF,12'h7EF},
{12'h8EF,12'h9EF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hFFF,12'h8FF,12'h8EF,12'h7EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'h8DF,12'h8EF,12'h8EF,12'h7DF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8FF,12'h7EF,12'h8EF,12'hDFF,12'hDFF,12'hDFF,12'hEFF,12'hDFF,12'hCFF,12'hCFF,12'hDFF,12'hDFF,12'hDFF,12'hDFF,12'h7FF,12'hDFF,12'hDFF,12'hBEF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hCFF,12'hEFF,12'hEFF,12'hBFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'h8EF,12'h8EF,12'h8EF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hCFF,12'hDFF,12'hEFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hCFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'h7EF,12'h8FF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hCFF,12'hDFF,12'hEFF,12'hCFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'h8FF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'hDFF,12'hCFF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h7DF,12'hDFF,12'hBFF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hCFF,12'hDFF,12'hDFF,12'hDFF,12'hCFF,12'hBFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hDFF,12'hDFF,12'hDFF,12'hBFF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'hDFF,12'hDFF,12'hDFF,12'hCFF,12'hDFF,12'hDFF,12'hCFF,12'hEFF,12'hDFF,12'hDFF,12'hDFF,12'hCFF,12'hCFF,12'hCFF,12'hDFF,12'hCFF,12'hDFF,12'hDFF,12'hCFF,12'h9EF,12'h7DF,12'h7DF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h7DF,12'hBFF,12'hCFF,12'h8FF,12'h8FF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'hAFF,12'hDFF,12'hDFF,12'hCFF,12'hDFF,12'hDFF,12'hBFF,12'hBEF,12'h9EF,12'h8EF,12'h8FF,12'h9DF,12'h8EF,12'h8FF,12'h8FF,12'h8EF,12'h8FF,12'h8EF,12'h8FF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hDFF,12'hDFF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h9EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h9EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h9EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hEFF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h9FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hFFF,12'hFFF,12'h8EF,12'h8EF,12'h8EF,12'hAEF,12'hEFF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h9EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h8FF,12'h8DF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8DF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8EF,12'h8EF,12'h9FF,12'h9EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hAEF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'hBDF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'h9FF,12'h9FF,12'h9EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h9EF,12'h9FF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDFF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hFFF,12'hFFF,12'hEFF,12'h8EF,12'h9EF,12'hFFF,12'hFFF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h9FF,12'h8EF,12'h8EF,12'h8FF,12'h8EF,12'h8EF,12'h9DF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'h8FF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'h8FF,12'hACF,12'hFFF,12'h8EF,12'h9EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'h8EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hCEF,12'h8EF,12'hFFF,12'hFFF,12'h8EF,12'h8EF,12'hAEF,12'h8FF,12'h8EF,12'h8FF,12'h8FF,12'h8EF,12'h8EF,12'h8EF,12'h8EF},
{12'h9EF,12'h9EF,12'h9FF,12'h8FF,12'h9EF,12'h9FF,12'h9EF,12'hFFF,12'hFFF,12'h8EF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'h8EF,12'h8FF,12'h9EF,12'h8FF,12'h9EF,12'h9EF,12'h9FF,12'h8EF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h9FF,12'h8FF,12'h8EF,12'h8FF,12'h8FF,12'h9EF,12'h9EF,12'h9EF,12'h8FF,12'h9EF,12'h9EF,12'h8FF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'h9EF,12'h9FF,12'h8FF,12'h9FF,12'h9EF},
{12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'hFFF,12'hBDF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'h8EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'h8EF,12'h9EF,12'h9FF,12'h9FF,12'h9FF},
{12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'h9EF,12'h9FF,12'h9EF,12'h9FF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hAEF,12'h9DF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'h9EF,12'h9FF,12'h9EF},
{12'h9FF,12'h9EF,12'h9EF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hCFF,12'hEFF,12'hEFF,12'hBFF,12'hEFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hDFF,12'hDFF,12'hDFF,12'hAEF,12'h9EF,12'h9FF,12'h9FF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'h9FF,12'h9FF,12'h9FF,12'hADF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'h9EF,12'h9EF,12'h9FF},
{12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h8EF,12'h8EF,12'hDEF,12'hCFF,12'hDFF,12'hDFF,12'hEFF,12'hCFF,12'hBEF,12'hCFF,12'hDFF,12'hCFF,12'hBFF,12'hCFF,12'hCFF,12'hBFF,12'hDFF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'hDFF,12'hDFF,12'hDFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hDFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hCFF,12'hDFF,12'hCFF,12'hDFF,12'hCFF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'hAEF,12'hBFF,12'hBEF,12'hDFF,12'hDFF,12'hDFF,12'hCFF,12'hDFF,12'hDFF,12'hDFF,12'hDFF,12'h9EF,12'h8EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF},
{12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'hCFF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h8EF,12'h9FF,12'h9EF,12'h9EF,12'hDFF,12'hDFF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9EF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF},
{12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF},
{12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF},
{12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'hAFF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'hAEF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF},
{12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'hAFF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF},
{12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF},
{12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'hFFF,12'hFFF,12'hAFF,12'h8EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'hAFF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'hAFF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'hAEF,12'h9FF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9EF,12'h9FF,12'h9EF,12'h9EF,12'h9EF,12'h9EF},
{12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hAFF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'hAEF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'hFFF,12'hFFF,12'hFFF,12'hDFF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'hFFF,12'hFFF,12'hFFF,12'h9EF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF,12'h9FF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'h9FF,12'hFFF,12'hFFF,12'h9EF,12'hAFF,12'hAFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h9FF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'h9FF,12'h9FF,12'h9EF,12'hAFF,12'h9FF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'h9FF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'h9FF,12'hAFF,12'hAFF,12'hAFF,12'h9FF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'h9FF,12'hFFF,12'hADF,12'hAFF,12'h9FF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'h9FF,12'hAFF,12'hAFF,12'h9EF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'h9FF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'h9FF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'h9FF,12'hAFF,12'hAFF,12'h9FF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'h9FF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hAEF,12'h9FF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hAFF,12'hAFF,12'hAEF,12'hFFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hAFF,12'hAEF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hCEF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBEF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'h9EF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'h9EF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'h9EF,12'hFFF,12'hAEF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFEF,12'hCFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'h9EF,12'hEFF,12'hEFF,12'hDFF,12'hBEF,12'hDFF,12'hDFF,12'hEFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hCFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hCEF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hDFF,12'hDFF,12'hDFF,12'hCEF,12'hCFF,12'hEFF,12'hEFF,12'hCFF,12'hDFF,12'hCFF,12'hEFF,12'hCFF,12'hCFF,12'hCEF,12'hBFF,12'h9EF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hAEF,12'hAFF,12'hAFF,12'hAFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hDFF,12'hDFF,12'hEFF,12'hDFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hDFF,12'hDFF,12'hEFF,12'hDFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hAFF,12'hAFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hCFF,12'hBFF,12'hAEF,12'hDFF,12'hDFF,12'hCFF,12'hBFF,12'hDFF,12'hDFF,12'hCFF,12'hBFF,12'hDFF,12'hBEF,12'hDFF,12'hDFF,12'hDFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hDFF,12'hDFF,12'hDFF,12'hDFF,12'hAEF,12'hDFF,12'hAFF,12'hCFF,12'hDFF,12'hDFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAEF,12'hAEF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hFFF,12'hFFF,12'hBDF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF},
{12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hAEF,12'hFFF,12'hFFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hDFF,12'hFFF,12'hFFF,12'hAFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hBFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hFFF,12'hAEF,12'hBEF,12'hFFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hBFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hBFF,12'hFFF,12'hCEF,12'hBFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hAFF,12'hAFF,12'hAFF,12'hBFF,12'hAFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hAEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hFFF,12'hBEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hBFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hAEF,12'hBFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBEF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hBEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hBEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hAEF,12'hFFF,12'hFFF,12'hBFF,12'hAEF,12'hFFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hADF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hEFF,12'hEFF,12'hEFF,12'hCFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hEFF,12'hEFF,12'hCFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hAFF,12'hAEF,12'hBFF,12'hBFF,12'hBFF,12'hAFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hAFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hEFF,12'hAEF,12'hFFF,12'hBEF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hFFF,12'hEFF,12'hBFF,12'hEFF,12'hDFF,12'hBEF,12'hCFF,12'hDFF,12'hCFF,12'hEFF,12'hEFF,12'hEFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBEF,12'hCFF,12'hCFF,12'hBFF,12'hBFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hCFF,12'hBFF,12'hDFF,12'hDFF,12'hDFF,12'hDFF,12'hBFF,12'hCFF,12'hCFF,12'hBFF,12'hEFF,12'hBFF,12'hBFF,12'hBFF,12'hDFF,12'hEFF,12'hEFF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hCFF,12'hAEF,12'hAEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hDFF,12'hBFF,12'hEFF,12'hEFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hDFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hBFF,12'hFFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hBEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hDFF,12'hEFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBEF,12'hEFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hBFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hEFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hCEF,12'hBEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hFFF,12'hDFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hBEF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hBEF,12'hBFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hCEF,12'hFFF,12'hEFF,12'hFFF,12'hFFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hBFF,12'hBFF,12'hBEF,12'hFFF,12'hFFF,12'hEFF,12'hEFF,12'hFFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hBDF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hEFF,12'hBFF,12'hBFF,12'hCFF,12'hBFF,12'hBEF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hFFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hCEF,12'hEFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hFFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hBFF,12'hBDF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hBEF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hCFF,12'hCFF,12'hCFF,12'hBEF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hFFF,12'hBFF,12'hBFF,12'hFFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hEFF,12'hCFF,12'hBFF,12'hCFF,12'hBEF,12'hDFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hEFF,12'hEFF,12'hEFF,12'hDFF,12'hDFF,12'hBFF,12'hBFF,12'hBFF,12'hBEF,12'hBFF,12'hCFF,12'hCEF,12'hDFF,12'hDFF,12'hDFF,12'hDFF,12'hCEF,12'hBFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hDFF,12'hDFF,12'hDFF,12'hDFF,12'hDFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hBFF},
{12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hBEF,12'hBFF,12'hDFF,12'hCFF,12'hDFF,12'hDFF,12'hBFF,12'hBFF,12'hBFF,12'hCFF,12'hCEF,12'hDFF,12'hCFF,12'hBFF,12'hBFF,12'hCFF,12'hDFF,12'hBFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hDFF,12'hDFF,12'hCFF,12'hCFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF,12'hBFF},
{12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hBFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hBFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF},
{12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hBFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF},
{12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF},
{12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF},
{12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF,12'hCFF}};
always @(posedge clk) begin
		if (pxl_y<80) begin
			background_drawing<=1;
			Red_background<=4'h7;
			Green_background<=4'hE;
			Blue_background <=4'hF;
		end
		else if (pxl_y>=80 && pxl_y<240) begin
			background_drawing<=1;
			Red_background <= Bitmap[{pxl_y}%80][{pxl_x}%80] [11:8];
			Green_background <= Bitmap[{pxl_y}%80][{pxl_x}%80] [7:4];
			Blue_background <= Bitmap[{pxl_y}%80][{pxl_x}%80] [3:0];
			

		end
			
		else begin 
		
			background_drawing<=1;
			Red_background<=4'hC;
			Green_background<=4'hF;
			Blue_background<=4'hF;
			
		end
		
			
		
			

end
endmodule
